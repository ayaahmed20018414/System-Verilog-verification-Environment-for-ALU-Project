//package includes files to be import easy
package ALU_pkg;
`include "transaction.svh"
`include "generator.svh"
`include "driver.svh"
`include "monitor.svh"
`include "scoreboard.svh"
`include "coverpoints.svh"
endpackage 
